TITLE
+ TITLE CONTINUES>...?
C1 3 6 1pF
R2 6 
   + 3 1k
.DC
;asdfasdfa
R5 +1 6 6;
*R5 1 6 3


*R5 1 6 6;
+FOOFLY

SUBCKT as asdf
R1 1 1 1 1  1
R2 3 43 34 3 3 
.ENDS


SUBCKT
.ENDS

.END

C1 1 1 1 