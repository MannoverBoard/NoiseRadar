Directive errors

C1 3 6 1pF


SUBCKT as asdf
SUBCKT
.ENDS
.ENDS

UNKNOWN DIRECTIVE


.ENDS

SUBCKT


.END

C1 1 1 1 1

